LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.std_logic_UNSIGNED.ALL;

ENTITY SR_REG IS
	PORT (		SET		: 				IN STD_LOGIC; 
				RESET	: 				IN STD_LOGIC;  
				OUTPUT	: 				OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE behavioral OF SR_REG IS

BEGIN
	PROCESS(SET, RESET)
	BEGIN
		IF(SET = '1'AND SET'EVENT)THEN
			OUTPUT <= '1';
		ELSIF (RESET = '1' AND RESET'EVENT) THEN
			OUTPUT <= '0';
		END IF;
		
	END PROCESS;
END behavioral;

