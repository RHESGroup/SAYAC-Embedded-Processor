module fulladder(i0, i1, ci, s, co);

wire S0;
wire S1;
wire S2;
wire S3;
wire S4;
wire S5;
wire S6;
wire S7;
wire S8;
wire S9;
wire S10;
wire S11;
wire S12;
wire S13;
wire S14;
wire S15;
wire S16;
input i0;
input i1;
input ci;
output s;
output co;

nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_0_ (
  .in1({ S12, S15 }),
  .out1({ S11 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1_ (
  .in1({ S10, S8 }),
  .out1({ S0 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2_ (
  .in1({ S12, S15 }),
  .out1({ S1 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3_ (
  .in1({ S1 }),
  .out1({ S2 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4_ (
  .in1({ S2, S11 }),
  .out1({ S3 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5_ (
  .in1({ S1, S0 }),
  .out1({ S4 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6_ (
  .in1({ S4, S14 }),
  .out1({ S5 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_7_ (
  .in1({ S3, S9 }),
  .out1({ S6 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_8_ (
  .in1({ S6, S5 }),
  .out1({ S16 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_9_ (
  .in1({ S0, S14 }),
  .out1({ S7 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_10_ (
  .in1({ S7, S1 }),
  .out1({ S13 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_11_ (
  .in1({ S15 }),
  .out1({ S8 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_12_ (
  .in1({ S14 }),
  .out1({ S9 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_13_ (
  .in1({ S12 }),
  .out1({ S10 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_14_ (
  .in1({ ci }),
  .out1({ S12 })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_15_ (
  .in1({ S13 }),
  .out1({ co })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_16_ (
  .in1({ i0 }),
  .out1({ S14 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_17_ (
  .in1({ i1 }),
  .out1({ S15 })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_18_ (
  .in1({ S16 }),
  .out1({ s })
);

endmodule