LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.std_logic_UNSIGNED.ALL;

ENTITY PARITY_GENERATOR IS
	GENERIC(	len					: INTEGER := 8);
	PORT (		DATA				: IN STD_LOGIC_VECTOR(len-1 downto 0);
				DATA_LEN_FORPARITY	: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
				PARITI_EVENODD		: IN STD_LOGIC;	
				PARITY				: OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE behavioral OF PARITY_GENERATOR IS
SIGNAL XOR_OUT : STD_LOGIC;



BEGIN
PARITY_PROCESS:	PROCESS (DATA, PARITI_EVENODD, DATA_LEN_FORPARITY)
BEGIN
	IF ( DATA_LEN_FORPARITY = "0101") THEN
		XOR_OUT <= DATA(0) XOR DATA(1) XOR DATA(2) XOR DATA(3) XOR DATA(4);
	ELSIF (DATA_LEN_FORPARITY = "0110")THEN
		XOR_OUT <= DATA(0) XOR DATA(1) XOR DATA(2) XOR DATA(3) XOR DATA(4) XOR DATA(5);
	ELSIF (DATA_LEN_FORPARITY = "0111")THEN
		XOR_OUT <= DATA(0) XOR DATA(1) XOR DATA(2) XOR DATA(3) XOR DATA(4) XOR DATA(5) XOR DATA(6);
	ELSIF (DATA_LEN_FORPARITY = "1000")THEN
		XOR_OUT <= DATA(0) XOR DATA(1) XOR DATA(2) XOR DATA(3) XOR DATA(4) XOR DATA(5)XOR DATA(6) XOR DATA(7);
	END IF;
	
	IF (PARITI_EVENODD = '1') THEN --EVEN PARITY
		IF (XOR_OUT = '1') THEN
			PARITY <= '1';
		ELSE PARITY <= '0';
		END IF;
	
	ELSIF (PARITI_EVENODD = '0') THEN --ODD PARITY
		IF (XOR_OUT = '1') THEN
			PARITY <= '0';
		ELSE PARITY <= '1';	
		END IF;
		
	END IF;
END PROCESS PARITY_PROCESS;
			
END behavioral;

