LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
 
ENTITY TB_PPI IS
	GENERIC( len		: INTEGER := 8;
			 len_bit	: INTEGER := 1);
END ENTITY;
 
ARCHITECTURE behavieral of TB_PPI is
    
   
SIGNAL CLK      : std_logic := '0';
SIGNAL rst      : std_logic := '0';
SIGNAL nRD		: STD_LOGIC; --READ SIGNAL
SIGNAL nWR		: STD_LOGIC; --WRITE SIGNAL
SIGNAL nCS		: STD_LOGIC; --CHIP SELECT
SIGNAL A		: std_logic_vector (1 downto 0); --PORT ADDRESS
SIGNAL PD		: std_logic_vector (len-1 downto 0); --PORT D
SIGNAL PA		: std_logic_vector (len-1 downto 0); --PORT A
SIGNAL PB		: std_logic_vector (len-1 downto 0); --PORT B
SIGNAL PCL		: std_logic_vector ((len/2)-1 downto 0); --PORTC LSB
SIGNAL PCU		: std_logic_vector ((len/2)-1 downto 0);
SIGNAL FLAG_TEST:  STD_LOGIC;

BEGIN

PPI_T1:ENTITY WORK.PPI2
	GENERIC MAP(len, len_bit	)
	PORT MAP(CLK, rst, nRD, nWR, nCS, A, PD, PA, PB, PCL, PCU);
---------------------------------------------------------------------------
-------------------------BSR TESTING---------------------------------------
PROCESS
BEGIN
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nCS <= '0';
	rst <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	rst <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	--rst <= '0';
	--PD(7) <= '0';
	--PD(3 DOWNTO 1) <= "000";
	--PD(0) <= '1';
	--PD(6 DOWNTO 4) <= "000";
	--WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	--PD(0) <= '0';
	--WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	--PD(3 DOWNTO 1) <= "001";
	--PD(0) <= '1';
	--PD(6 DOWNTO 4) <= "000";
	--WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	--PD(0) <= '0';
	--WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	--PD(3 DOWNTO 1) <= "011";
	--PD(0) <= '1';
	--PD(6 DOWNTO 4) <= "000";
	--WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	--PD(0) <= '0';
---------------------------------------------------------------------------
-------------------------MODE0 TESTING-------------------------------------

	A <= "11"; --CONTROL REGISTER MODE
	PD <= "10010000"; ----GROUPA SIMPLE I/O (PA IS INPUT)
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PD <= (OTHERS => 'Z');
	A <= "00";
	PA <= "11110111";
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '1';
	PA <= (OTHERS => 'Z');
	
	A <= "11"; --CONTROL REGISTER MODE
	PD <= "10000000"; ----GROUPA SIMPLE I/O (PA IS OUTPUT)
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PD <= (OTHERS => 'Z');
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PD <= "10101010";
	A <= "00";
	nWR <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nWR <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nWR <= '1';
	
	A <= "11"; --CONTROL REGISTER MODE
	PD <= "10001000"; ----GROUPA SIMPLE I/O (PCU IS INPUT)
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PD <= (OTHERS => 'Z');
	A <= "10";
	PCU <= "1001";
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '1';
	PCU <= (OTHERS => 'Z');
	
	A <= "11"; --CONTROL REGISTER MODE
	PD <= "10000000"; ----GROUPA SIMPLE I/O (PCU IS OUTPUT)
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PD <= (OTHERS => 'Z');
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PD <= "11110000";
	A <= "10";
	nWR <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nWR <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nWR <= '1';
	
	
	A <= "11"; --CONTROL REGISTER MODE
	PD <= "10000010"; ----GROUPB SIMPLE I/O (PB IS INPUT)
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PD <= (OTHERS => 'Z');
	A <= "01";
	PB <= "10011001";
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '1';
	PB <= (OTHERS => 'Z');
	
	A <= "11"; --CONTROL REGISTER MODE
	PD <= "10000000"; ----GROUPB SIMPLE I/O (PB IS OUTPUT)
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PD <= (OTHERS => 'Z');
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PD <= "10000001";
	A <= "01";
	nWR <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nWR <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nWR <= '1';
	
	A <= "11"; --CONTROL REGISTER MODE
	PD <= "10000001"; ----GROUPB SIMPLE I/O (PCL IS INPUT)
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PD <= (OTHERS => 'Z');
	A <= "10";
	PCL <= "1010";
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '1';
	PCL <= (OTHERS => 'Z');
	
	A <= "11"; --CONTROL REGISTER MODE
	PD <= "10000000"; ----GROUPB SIMPLE I/O (PCU IS OUTPUT)
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PD <= (OTHERS => 'Z');
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PD <= "10011101";
	A <= "10";
	nWR <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nWR <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nWR <= '1';
	PD <= (OTHERS => 'Z');
	A <="ZZ";
-------------------------------------------------------------------------
-----------------------MODE1 TESTING-------------------------------------	
	rst <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	rst <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	rst <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	A <= "11"; --CONTROL REGISTER MODE
	PD <= "10110000"; ----GROUPA STROBED I/O (PA IS INPUT)
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PD <= (OTHERS => 'Z');
	PA <= "10010000";
	A <= "ZZ";
	PCU(0) <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PCU(0) <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PCU(0) <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '1';
	
	PD <= (OTHERS => 'Z');
	PA <= (OTHERS => 'Z');
	PCU<= (OTHERS => 'Z');
	PCL <=(OTHERS => 'Z');
	rst <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	rst <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	rst <= '0';
	A <= "11"; --CONTROL REGISTER MODE
	PCU(2) <= '1';
	PD <= "10100000"; ----GROUPA STROBED I/O (PA IS OUTPUT)
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	A <= "ZZ";
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PD <="11100011";
	nWR <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nWR <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nWR <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PCU(2) <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PCU(2) <= '1';
	
	
	PD <= (OTHERS => 'Z');
	PA <= (OTHERS => 'Z');
	PCU<= (OTHERS => 'Z');
	PCL <=(OTHERS => 'Z');
	rst <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	rst <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	rst <= '0';
	A <= "11"; --CONTROL REGISTER MODE
	PD <= "10000110"; ----GROUPB STROBED I/O (PB IS INPUT)
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PD <= (OTHERS => 'Z');
	PB <= "10010000";
	A <= "ZZ";
	PCL(2) <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PCL(2) <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PCL(2) <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '1';
	
	PD <= (OTHERS => 'Z');
	PA <= (OTHERS => 'Z');
	PCU<= (OTHERS => 'Z');
	PCL <=(OTHERS => 'Z');
	PB <=(OTHERS => 'Z');
	rst <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	rst <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	rst <= '0';
	A <= "11"; --CONTROL REGISTER MODE
	PD <= "10000100"; ----GROUPA STROBED I/O (PB IS OUTPUT)
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PCL(2) <= '1';
	A <= "ZZ";
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PD <="11001100";
	nWR <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nWR <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nWR <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PCL(2) <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PCL(2) <= '1';
	
---------------------------------------------------------------------------
-------------------------MODE2 TESTING-------------------------------------	
	PD <= (OTHERS => 'Z');
	PA <= (OTHERS => 'Z');
	PCU<= (OTHERS => 'Z');
	PCL <=(OTHERS => 'Z');
	PB <=(OTHERS => 'Z');
	rst <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	rst <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	rst <= '0';
	A <= "11"; --CONTROL REGISTER MODE
	PD <= "11010000"; ----GROUPA BIDIRECTIONAL I/O(INPUT OPERATION)
	PCU(0) <= '1';
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	A <= "ZZ";
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PA <="11110000";
	PCU(0)<= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PCU(0)<= '1';
	
	PD <= (OTHERS => 'Z');
	PA <= (OTHERS => 'Z');
	PCU<= (OTHERS => 'Z');
	PCL <=(OTHERS => 'Z');
	PB <=(OTHERS => 'Z');
	rst <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	rst <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	rst <= '0';
	A <= "11"; --CONTROL REGISTER MODE
	PD <= "11000000"; ----GROUPA BIDIRECTIONAL I/O(OUTPUT OPERATION)
	PCU(2) <= '1';
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nRD <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	A <= "ZZ";
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PD <="11110111";
	nWR <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nWR <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	nWR <= '1';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PCU(2) <= '0';
	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);	WAIT UNTIL (CLK = '1' AND CLK'EVENT); WAIT UNTIL (CLK = '1' AND CLK'EVENT);
	PCU(2) <= '0';
	WAIT FOR 1000 ns;
END PROCESS;
--------------------------------------------------------------------------	
setclk: PROCESS
		BEGIN
			WAIT FOR 5 NS;
			CLK <= NOT clk;
			WAIT FOR 5 NS;
		END PROCESS setclk;
END behavieral;