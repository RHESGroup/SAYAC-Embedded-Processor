LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
 
ENTITY TB_UART2 IS
	GENERIC( COUNTER_RANGE	:	INTEGER	:=	87;
			 len			:	INTEGER	:=	8;
			 Cnt_len		:	INTEGER	:=	4;
			 DATA_SERIAL_len:	INTEGER	:=	8);
END ENTITY;
 
ARCHITECTURE behavieral of TB_UART2 is
    
  -- Test Bench uses a 10 MHz Clock
  -- Want to interface to 115200 baud UART
  -- 10000000 / 115200 = 87 Clocks Per Bit.
SIGNAL CLK   :   STD_LOGIC:= '0';    			
SIGNAL rst   :   STD_LOGIC;
SIGNAL nWR   :   STD_LOGIC;
SIGNAL nRD   :   STD_LOGIC;
SIGNAL CD    :   STD_LOGIC;
SIGNAL nCS   :   STD_LOGIC;
SIGNAL nCTS  :   STD_LOGIC; --ACTIVE LOW CLEAAR TO SEND SERIAL DATA
SIGNAL DATA  : 	 STD_LOGIC_VECTOR(len-1 downto 0); --r_TX_BYTE / w_RX_BYTE
SIGNAL TXE   :   STD_LOGIC; --TRANSMITTER EMPTY
SIGNAL TXRDY :   STD_LOGIC; --TRANSMITTER EMPTY
SIGNAL RXRDY :   STD_LOGIC; --TRANSMITTER EMPTY
SIGNAL TXD 	 :   STD_LOGIC; --DATA SERIAL TRANSFER
SIGNAL BREAK :   STD_LOGIC; --GOES HIGH WHEN HAVE 2 STOP BIT 
SIGNAL DATA_LEN_FORPARITY	: STD_LOGIC_VECTOR(3 DOWNTO 0);        
SIGNAL PARITI_EVENODD		: STD_LOGIC;	
SIGNAL PARITY				: STD_LOGIC;
BEGIN
	
CLK <= not CLK after 50 ns;
 
CHIP_INST:ENTITY WORK.CHIP 
	GENERIC MAP( COUNTER_RANGE, len, Cnt_len, DATA_SERIAL_len)
	PORT MAP(CLK, rst, nWR, nRD, CD, nCS, nCTS, DATA , TXE , TXRDY, RXRDY, BREAK);	
	
--PARITY_INST:ENTITY WORK.PARITY_GENERATOR 
--	GENERIC MAP(len)
--	PORT MAP(DATA, DATA_LEN_FORPARITY, PARITI_EVENODD, PARITY);	
--TEST_PARITY: PROCESS
--BEGIN
--
--DATA <= "10101010";
--DATA_LEN_FORPARITY <= "1000";
--PARITI_EVENODD <= '0';
--
--WAIT FOR 100 NS;
--
--END PROCESS TEST_PARITY;
--TX_INST: entity WORK.UART_TX 
--  GENERIC MAP(COUNTER_RANGE,  len,	Cnt_len)
--  PORT MAP(Clk, rst, nCS, nCTS, CD, nWR, DATA, TXD, TXE );



TEST_TX: PROCESS
BEGIN
nCS <= '0';
WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);
nWR <= '1';
CD <= '1';
DATA <= "01010010";
WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);
nWR <= '0';	
WAIT UNTIL (CLK = '1' AND CLK'EVENT);
nWR <= '1';	
CD <= '0';
DATA <= "10101011";
WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);
nWR <= '0';	
WAIT UNTIL (CLK = '1' AND CLK'EVENT);
nWR <= '1';
WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);
nCTS <= '0';
WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);
DATA <= (OTHERS => 'Z');
nRD <= '1';
WAIT UNTIL (CLK = '1' AND CLK'EVENT);WAIT UNTIL (CLK = '1' AND CLK'EVENT);
nRD <= '0';
WAIT FOR 10000000 NS;
END PROCESS TEST_TX;


	  
end behavieral;
