LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
 
ENTITY TB_COUNTER IS
	GENERIC( LEN_CONTROLWORD	: INTEGER := 6;
			 LEN_DATA			: INTEGER := 8;
			 len				: INTEGER := 16);
END ENTITY;
 
ARCHITECTURE behavieral of TB_COUNTER is
    
   
SIGNAL CLK_INPUT			: STD_LOGIC := '0';
SIGNAL rst					: STD_LOGIC;
SIGNAL CONTROLWORD			: STD_LOGIC_VECTOR (5 DOWNTO 0);
SIGNAL GATE					: STD_LOGIC;
SIGNAL WR_SIGNAL			: STD_LOGIC;
SIGNAL RD_SIGNAL			: STD_LOGIC;
SIGNAL STATUS_RD			: STD_LOGIC;--ENABLESTATUSLATCH
SIGNAL RD_BACK				: STD_LOGIC;--EnableCounterLatch
SIGNAL DATABUS				: STD_LOGIC_VECTOR (LEN_DATA-1 DOWNTO 0);
SIGNAL OUTPUT				: STD_LOGIC;
SIGNAL NUM_IN				: STD_LOGIC_VECTOR(len-1 downto 0);
SIGNAL DOWN_COUNT_BINARY	: STD_LOGIC;
SIGNAL DOWN_COUNT_BCD		: STD_LOGIC;
SIGNAL LOAD_NUMIN			: STD_LOGIC;
SIGNAL MODE					: STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL FLAGOUT_DURATION		: STD_LOGIC;
SIGNAL NUM_OUT				: STD_LOGIC_VECTOR(len-1 downto 0);
SIGNAL DATA					: STD_LOGIC_VECTOR(LEN_DATA-1 downto 0);
SIGNAL RD					: STD_LOGIC;
SIGNAL WR					: STD_LOGIC;
SIGNAL CS					: STD_LOGIC;
SIGNAL A0					: STD_LOGIC;
SIGNAL A1					: STD_LOGIC;
SIGNAL GATE0				: STD_LOGIC;
SIGNAL GATE1				: STD_LOGIC;
SIGNAL GATE2				: STD_LOGIC;
SIGNAL OUT0					: STD_LOGIC;
SIGNAL OUT1					: STD_LOGIC;
SIGNAL OUT2					: STD_LOGIC;

BEGIN

CHIP_INST:ENTITY WORK.CHIP
	GENERIC MAP(LEN_CONTROLWORD, LEN_DATA)
	PORT MAP(DATA, RD, WR, CS, A0, A1, CLK_INPUT, CLK_INPUT, CLK_INPUT,	rst, GATE0,	GATE1, GATE2, OUT0,	OUT1, OUT2);
	
-------------------------------------------------------------------------------------
--------------------------------CHIP TESTING-----------------------------------------
PROCESS
BEGIN

WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
rst <= '0';
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT); WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
rst <= '1';
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT); WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
rst <= '0';
CS <= '1';
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
CS <= '0';
A1 <= '1'; A0 <= '1';
WR <= '0'; RD <= '1';
DATA <= "00111010";
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
WR <= '1'; RD <= '1';
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
WR <= '0'; RD <= '1';
A1 <= '0'; A0 <= '0';
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
WR <= '1'; RD <= '1';
DATA <= "00001111";
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
DATA <= "00000000";
GATE0 <= '0';
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
GATE0 <= '1';
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND 
CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
GATE0 <= '0';
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
GATE0 <= '1';
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);

WR <= '0'; RD <= '1';
A1 <= '0'; A0 <= '0';
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
WR <= '1'; RD <= '1';
DATA <= "00000111";
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
DATA <= "00000000";
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
DATA <= (OTHERS => 'Z');
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);


A1 <= '1'; A0 <= '1';
WR <= '0'; RD <= '1';
DATA <= "11110011";
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
WR <= '1'; RD <= '1';
DATA <= (OTHERS => 'Z');
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
A1 <= '0'; A0 <= '0';
WR <= '1'; RD <= '0';
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
WR <= '1'; RD <= '1';
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
A1 <= '1'; A0 <= '1';
WR <= '0'; RD <= '1';
DATA <= "11000011";
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
DATA <= (OTHERS => 'Z');
WR <= '1'; RD <= '1';
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
A1 <= '0'; A0 <= '0';
WR <= '1'; RD <= '0';
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
WR <= '1'; RD <= '1';
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
WR <= '1'; RD <= '0';
WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
WR <= '1'; RD <= '1';
DATA <= (OTHERS => 'Z');


WAIT FOR 1000 ns;
END PROCESS;

--------------------------------------------------------------------------------------		
	
--Counter_T1:ENTITY WORK.Counter
--	GENERIC MAP( LEN_CONTROLWORD, LEN_DATA)
--	PORT MAP(CLK_INPUT, rst	, CONTROLWORD, GATE	, WR_SIGNAL	, RD_SIGNAL	, STATUS_RD	, RD_BACK, DATABUS, OUTPUT);
	
-------------------------------------------------------------------------
-------------------------TESTING COUNTER---------------------------------------
--PROCESS
--BEGIN
--	WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT); WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT); WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
--	rst <= '0';
--	WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT); WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
--	rst <= '1';
--	WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT); WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
--	rst <= '0';
--	--GATE <= '0';
--	WR_SIGNAL <= '0';
--	CONTROLWORD <= "110011"; --LSB ONLY MODE0 BINARY
--	--DATABUS <= "00001111";
--	WR_SIGNAL <= '0';
--	WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
--	WR_SIGNAL <= '1';
--	WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
--	WR_SIGNAL <= '0';
--	DATABUS <= "00000111";
--	WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
--	DATABUS <= "00000000";
--	WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
--	--WR_SIGNAL <= '1';
--	--WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
--	WR_SIGNAL <= '0';
--	--DATABUS <= "11000111";
--	WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
--	--DATABUS <= "00000000";
--	GATE <= '1';
--	WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
--	--GATE <= '1';
--	WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
--	--GATE <= '0';
--	WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
--	--GATE <= '1';
--	WR_SIGNAL <= '1';
--	WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
--	WR_SIGNAL <= '0';
--	DATABUS <= "00001111";
--	WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
--	DATABUS <= "00000000";
--	WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
--	GATE <= '0';
--	WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
--	
--	--GATE <= '1';
--	WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
--	--GATE <= '0';
--	WAIT FOR 1000 ns;
--END PROCESS;
----------------------------------------------------------------------------------------
-----------------------------DOWN_COUNTER TESTING---------------------------------------
--DOWN_COUNTER_INST:ENTITY WORK.DOWN_COUNTER 
--	GENERIC MAP(len)
--	PORT MAP(CLK_INPUT, rst, NUM_IN, DOWN_COUNT_BINARY, DOWN_COUNT_BCD, LOAD_NUMIN, MODE, FLAGOUT_DURATION, NUM_OUT);
----DOWN_COUNTER_TEST: PROCESS
--BEGIN
--	NUM_IN <= "0000000000000111";
--	MODE <= "000";
--	WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
--	LOAD_NUMIN <= '1';
--	WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
--	LOAD_NUMIN <= '0';
--	WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
--	DOWN_COUNT_BINARY <= '1';
--	WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
--	DOWN_COUNT_BINARY <= '0';
--	WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
--	DOWN_COUNT_BINARY <= '1';
--	WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
--	DOWN_COUNT_BINARY <= '0';
--	WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
--	DOWN_COUNT_BINARY <= '1';
--	WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
--	DOWN_COUNT_BINARY <= '0';
--	WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
--	DOWN_COUNT_BINARY <= '1';
--	WAIT UNTIL (CLK_INPUT = '1' AND CLK_INPUT'EVENT);
--	DOWN_COUNT_BINARY <= '0';
--	
--	
--	
--	WAIT FOR 1000 ns;
--END PROCESS;
-------------------------------------------------------------------------------------
--------------------------------CHIP TESTING-----------------------------------------
PROCESS
BEGIN



WAIT FOR 1000 ns;
END PROCESS;








--------------------------------------------------------------------------------------













	
setCLK_INPUT: PROCESS
		BEGIN
			WAIT FOR 5 NS;
			CLK_INPUT <= NOT CLK_INPUT;
			WAIT FOR 5 NS;
		END PROCESS setCLK_INPUT;
END behavieral;